module mult(in, out);

	input signed [8:0] in;
	parameter mult_num = 11'd1638;
	
	output signed [19:0] out;
	
	wire [8:0] in;
	wire [19:0] out;
	
	assign out = mult_num * in;

endmodule 